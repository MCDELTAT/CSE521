`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   10:44:40 01/18/2017
// Design Name:   bi_directional_shift
// Module Name:   /home/aaron/Git Repos/CSE311/lab1/bi_directional_shift_tb.v
// Project Name:  lab1
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: bi_directional_shift
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module bi_directional_shift_tb;

	// Inputs
	reg [7:0] d_in;
	reg [2:0] shift_amount;
	reg shift_direction;

	// Outputs
	wire [7:0] shifter_out;

	// Instantiate the Unit Under Test (UUT)
	bi_directional_shift uut (
		.d_in(d_in), 
		.shift_amount(shift_amount), 
		.shift_direction(shift_direction), 
		.shifter_out(shifter_out)
	);

	initial begin
		// Initialize Inputs
		d_in = 0;
		shift_amount = 0;
		shift_direction = 0;

		// Wait 100 ns for global reset to finish
		#100;
        
		// Test shift left 2
		shift_direction = 1'b0;
		d_in = 8'b00100000;
		shift_amount = 3'b010;
		
		#100;
		// Test shift right 3
		shift_direction = 1'b1;
		d_in = 8'b00010000;
		shift_amount = 3'b011;

	end
      
endmodule

